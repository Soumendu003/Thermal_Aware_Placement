--
--  Copyright (c) 2003 Launchbird Design Systems, Inc.
--  All rights reserved.
--  
--  Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
--    Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
--    Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
--  
--  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES,
--  INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED.
--  IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY,
--  OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
--  OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
--  (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
--  
--  
--  Overview:
--  
--    Low-density parity-check (LDPC) codes are forward error correction codes invented
--    by Robert Gallager in the early 60's.  Like turbo codes, LDPC codes approach Shannon's
--    limit for channel capacity, but have reduced decoding complexity.
--  
--  Architecture:
--  
--    This LDPC error corrector implements Gallager's "A" algorithm: an iterative,
--    hard-decision decoder that opts for simplicity over performance.  The architecture
--    elaborates all logic required to implement the message-passing algorithm from
--    message nodes, to check nodes, then back to message nodes -- one iteration occurs
--    every clock cycle.
--  
--    The core is primarily meant as an LDPC evaluation platform, as the fully parallel
--    architecture may be inappropriate for synthesizing large block length LDPC decoders.
--  
--    The LDPC code is defined by a parity check matrix, and is specified from the Confluence source.
--    This LDPC corrector has been generated for the following parity check matrix:
--  
--  1 1 1 1 . . . . . . . . . . . . . . . . 
--  . . . . 1 1 1 1 . . . . . . . . . . . . 
--  . . . . . . . . 1 1 1 1 . . . . . . . . 
--  . . . . . . . . . . . . 1 1 1 1 . . . . 
--  . . . . . . . . . . . . . . . . 1 1 1 1 
--  1 . . . 1 . . . 1 . . . 1 . . . . . . . 
--  . 1 . . . 1 . . . 1 . . . . . . 1 . . . 
--  . . 1 . . . 1 . . . . . . 1 . . . 1 . . 
--  . . . 1 . . . . . . 1 . . . 1 . . . 1 . 
--  . . . . . . . 1 . . . 1 . . . 1 . . . 1 
--  1 . . . . 1 . . . . . 1 . . . . . 1 . . 
--  . 1 . . . . 1 . . . 1 . . . . 1 . . . . 
--  . . 1 . . . . 1 . . . . 1 . . . . . 1 . 
--  . . . 1 . . . . 1 . . . . 1 . . 1 . . . 
--  . . . . 1 . . . . 1 . . . . 1 . . . . 1 
--  
--  
--  Interface:
--  
--    Synchronization:
--      clock_c      : Clock.
--  
--    Inputs:
--      start_i      : Start signal pulse.  Aligned with input message.
--      message_i    : Input message.
--  
--    Outputs:
--      valid_o      : High if output message meets parity checking.
--      message_o    : Output message.
--  
--  
--  
--  
--  
--  Generated by Confluence 0.6.3  --  Launchbird Design Systems, Inc.  --  www.launchbird.com
--  
--  Build Date : Fri Aug 22 09:48:55 CDT 2003
--  
--  Interface
--  
--    Build Name    : cf_ldpc
--    Clock Domains : clock_c  
--    Vector Input  : start_i(1)
--    Vector Input  : message_i(20)
--    Vector Output : valid_o(1)
--    Vector Output : message_o(20)
--  
--  
--  

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_103 is
port (
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(1 downto 0);
i3 : in  unsigned(1 downto 0);
o1 : out unsigned(1 downto 0));
end entity cf_ldpc_103;
architecture rtl of cf_ldpc_103 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(1 downto 0);
begin
n1 <= i1(1 downto 1);
n2 <= i2(1 downto 1);
n3 <= i3(1 downto 1);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(0 downto 0);
n6 <= i2(0 downto 0);
n7 <= i3(0 downto 0);
n8 <= n5(0 downto 0);
n9 <= n6(0 downto 0);
n10 <= n7(0 downto 0);
n11 <= n9 when n8 = "1" else n10;
n12 <= n4 & n11;
o1 <= n12;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_102 is
port (
i1 : in  unsigned(2 downto 0);
i2 : in  unsigned(2 downto 0);
i3 : in  unsigned(2 downto 0);
o1 : out unsigned(2 downto 0));
end entity cf_ldpc_102;
architecture rtl of cf_ldpc_102 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(1 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(1 downto 0);
signal n8 : unsigned(2 downto 0);
signal s9_1 : unsigned(1 downto 0);
component cf_ldpc_103 is
port (
i1 : in  unsigned(1 downto 0);
i2 : in  unsigned(1 downto 0);
i3 : in  unsigned(1 downto 0);
o1 : out unsigned(1 downto 0));
end component cf_ldpc_103;
begin
n1 <= i1(2 downto 2);
n2 <= i2(2 downto 2);
n3 <= i3(2 downto 2);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_103 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_101 is
port (
i1 : in  unsigned(3 downto 0);
i2 : in  unsigned(3 downto 0);
i3 : in  unsigned(3 downto 0);
o1 : out unsigned(3 downto 0));
end entity cf_ldpc_101;
architecture rtl of cf_ldpc_101 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(2 downto 0);
signal n6 : unsigned(2 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(3 downto 0);
signal s9_1 : unsigned(2 downto 0);
component cf_ldpc_102 is
port (
i1 : in  unsigned(2 downto 0);
i2 : in  unsigned(2 downto 0);
i3 : in  unsigned(2 downto 0);
o1 : out unsigned(2 downto 0));
end component cf_ldpc_102;
begin
n1 <= i1(3 downto 3);
n2 <= i2(3 downto 3);
n3 <= i3(3 downto 3);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_102 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_100 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(4 downto 0);
i3 : in  unsigned(4 downto 0);
o1 : out unsigned(4 downto 0));
end entity cf_ldpc_100;
architecture rtl of cf_ldpc_100 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(3 downto 0);
signal n6 : unsigned(3 downto 0);
signal n7 : unsigned(3 downto 0);
signal n8 : unsigned(4 downto 0);
signal s9_1 : unsigned(3 downto 0);
component cf_ldpc_101 is
port (
i1 : in  unsigned(3 downto 0);
i2 : in  unsigned(3 downto 0);
i3 : in  unsigned(3 downto 0);
o1 : out unsigned(3 downto 0));
end component cf_ldpc_101;
begin
n1 <= i1(4 downto 4);
n2 <= i2(4 downto 4);
n3 <= i3(4 downto 4);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_101 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_99 is
port (
i1 : in  unsigned(5 downto 0);
i2 : in  unsigned(5 downto 0);
i3 : in  unsigned(5 downto 0);
o1 : out unsigned(5 downto 0));
end entity cf_ldpc_99;
architecture rtl of cf_ldpc_99 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(4 downto 0);
signal n7 : unsigned(4 downto 0);
signal n8 : unsigned(5 downto 0);
signal s9_1 : unsigned(4 downto 0);
component cf_ldpc_100 is
port (
i1 : in  unsigned(4 downto 0);
i2 : in  unsigned(4 downto 0);
i3 : in  unsigned(4 downto 0);
o1 : out unsigned(4 downto 0));
end component cf_ldpc_100;
begin
n1 <= i1(5 downto 5);
n2 <= i2(5 downto 5);
n3 <= i3(5 downto 5);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_100 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_98 is
port (
i1 : in  unsigned(6 downto 0);
i2 : in  unsigned(6 downto 0);
i3 : in  unsigned(6 downto 0);
o1 : out unsigned(6 downto 0));
end entity cf_ldpc_98;
architecture rtl of cf_ldpc_98 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(5 downto 0);
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(5 downto 0);
signal n8 : unsigned(6 downto 0);
signal s9_1 : unsigned(5 downto 0);
component cf_ldpc_99 is
port (
i1 : in  unsigned(5 downto 0);
i2 : in  unsigned(5 downto 0);
i3 : in  unsigned(5 downto 0);
o1 : out unsigned(5 downto 0));
end component cf_ldpc_99;
begin
n1 <= i1(6 downto 6);
n2 <= i2(6 downto 6);
n3 <= i3(6 downto 6);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_99 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_97 is
port (
i1 : in  unsigned(7 downto 0);
i2 : in  unsigned(7 downto 0);
i3 : in  unsigned(7 downto 0);
o1 : out unsigned(7 downto 0));
end entity cf_ldpc_97;
architecture rtl of cf_ldpc_97 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(6 downto 0);
signal n6 : unsigned(6 downto 0);
signal n7 : unsigned(6 downto 0);
signal n8 : unsigned(7 downto 0);
signal s9_1 : unsigned(6 downto 0);
component cf_ldpc_98 is
port (
i1 : in  unsigned(6 downto 0);
i2 : in  unsigned(6 downto 0);
i3 : in  unsigned(6 downto 0);
o1 : out unsigned(6 downto 0));
end component cf_ldpc_98;
begin
n1 <= i1(7 downto 7);
n2 <= i2(7 downto 7);
n3 <= i3(7 downto 7);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_98 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_96 is
port (
i1 : in  unsigned(8 downto 0);
i2 : in  unsigned(8 downto 0);
i3 : in  unsigned(8 downto 0);
o1 : out unsigned(8 downto 0));
end entity cf_ldpc_96;
architecture rtl of cf_ldpc_96 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(7 downto 0);
signal n7 : unsigned(7 downto 0);
signal n8 : unsigned(8 downto 0);
signal s9_1 : unsigned(7 downto 0);
component cf_ldpc_97 is
port (
i1 : in  unsigned(7 downto 0);
i2 : in  unsigned(7 downto 0);
i3 : in  unsigned(7 downto 0);
o1 : out unsigned(7 downto 0));
end component cf_ldpc_97;
begin
n1 <= i1(8 downto 8);
n2 <= i2(8 downto 8);
n3 <= i3(8 downto 8);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_97 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_95 is
port (
i1 : in  unsigned(9 downto 0);
i2 : in  unsigned(9 downto 0);
i3 : in  unsigned(9 downto 0);
o1 : out unsigned(9 downto 0));
end entity cf_ldpc_95;
architecture rtl of cf_ldpc_95 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(8 downto 0);
signal n6 : unsigned(8 downto 0);
signal n7 : unsigned(8 downto 0);
signal n8 : unsigned(9 downto 0);
signal s9_1 : unsigned(8 downto 0);
component cf_ldpc_96 is
port (
i1 : in  unsigned(8 downto 0);
i2 : in  unsigned(8 downto 0);
i3 : in  unsigned(8 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_ldpc_96;
begin
n1 <= i1(9 downto 9);
n2 <= i2(9 downto 9);
n3 <= i3(9 downto 9);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_96 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_94 is
port (
i1 : in  unsigned(10 downto 0);
i2 : in  unsigned(10 downto 0);
i3 : in  unsigned(10 downto 0);
o1 : out unsigned(10 downto 0));
end entity cf_ldpc_94;
architecture rtl of cf_ldpc_94 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(9 downto 0);
signal n6 : unsigned(9 downto 0);
signal n7 : unsigned(9 downto 0);
signal n8 : unsigned(10 downto 0);
signal s9_1 : unsigned(9 downto 0);
component cf_ldpc_95 is
port (
i1 : in  unsigned(9 downto 0);
i2 : in  unsigned(9 downto 0);
i3 : in  unsigned(9 downto 0);
o1 : out unsigned(9 downto 0));
end component cf_ldpc_95;
begin
n1 <= i1(10 downto 10);
n2 <= i2(10 downto 10);
n3 <= i3(10 downto 10);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_95 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_93 is
port (
i1 : in  unsigned(11 downto 0);
i2 : in  unsigned(11 downto 0);
i3 : in  unsigned(11 downto 0);
o1 : out unsigned(11 downto 0));
end entity cf_ldpc_93;
architecture rtl of cf_ldpc_93 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(10 downto 0);
signal n6 : unsigned(10 downto 0);
signal n7 : unsigned(10 downto 0);
signal n8 : unsigned(11 downto 0);
signal s9_1 : unsigned(10 downto 0);
component cf_ldpc_94 is
port (
i1 : in  unsigned(10 downto 0);
i2 : in  unsigned(10 downto 0);
i3 : in  unsigned(10 downto 0);
o1 : out unsigned(10 downto 0));
end component cf_ldpc_94;
begin
n1 <= i1(11 downto 11);
n2 <= i2(11 downto 11);
n3 <= i3(11 downto 11);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_94 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_92 is
port (
i1 : in  unsigned(12 downto 0);
i2 : in  unsigned(12 downto 0);
i3 : in  unsigned(12 downto 0);
o1 : out unsigned(12 downto 0));
end entity cf_ldpc_92;
architecture rtl of cf_ldpc_92 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(11 downto 0);
signal n6 : unsigned(11 downto 0);
signal n7 : unsigned(11 downto 0);
signal n8 : unsigned(12 downto 0);
signal s9_1 : unsigned(11 downto 0);
component cf_ldpc_93 is
port (
i1 : in  unsigned(11 downto 0);
i2 : in  unsigned(11 downto 0);
i3 : in  unsigned(11 downto 0);
o1 : out unsigned(11 downto 0));
end component cf_ldpc_93;
begin
n1 <= i1(12 downto 12);
n2 <= i2(12 downto 12);
n3 <= i3(12 downto 12);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(11 downto 11) &
  i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_93 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_91 is
port (
i1 : in  unsigned(13 downto 0);
i2 : in  unsigned(13 downto 0);
i3 : in  unsigned(13 downto 0);
o1 : out unsigned(13 downto 0));
end entity cf_ldpc_91;
architecture rtl of cf_ldpc_91 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(12 downto 0);
signal n6 : unsigned(12 downto 0);
signal n7 : unsigned(12 downto 0);
signal n8 : unsigned(13 downto 0);
signal s9_1 : unsigned(12 downto 0);
component cf_ldpc_92 is
port (
i1 : in  unsigned(12 downto 0);
i2 : in  unsigned(12 downto 0);
i3 : in  unsigned(12 downto 0);
o1 : out unsigned(12 downto 0));
end component cf_ldpc_92;
begin
n1 <= i1(13 downto 13);
n2 <= i2(13 downto 13);
n3 <= i3(13 downto 13);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(12 downto 12) &
  i2(11 downto 11) &
  i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_92 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_90 is
port (
i1 : in  unsigned(14 downto 0);
i2 : in  unsigned(14 downto 0);
i3 : in  unsigned(14 downto 0);
o1 : out unsigned(14 downto 0));
end entity cf_ldpc_90;
architecture rtl of cf_ldpc_90 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(13 downto 0);
signal n6 : unsigned(13 downto 0);
signal n7 : unsigned(13 downto 0);
signal n8 : unsigned(14 downto 0);
signal s9_1 : unsigned(13 downto 0);
component cf_ldpc_91 is
port (
i1 : in  unsigned(13 downto 0);
i2 : in  unsigned(13 downto 0);
i3 : in  unsigned(13 downto 0);
o1 : out unsigned(13 downto 0));
end component cf_ldpc_91;
begin
n1 <= i1(14 downto 14);
n2 <= i2(14 downto 14);
n3 <= i3(14 downto 14);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(13 downto 13) &
  i2(12 downto 12) &
  i2(11 downto 11) &
  i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_91 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_89 is
port (
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_ldpc_89;
architecture rtl of cf_ldpc_89 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(14 downto 0);
signal n6 : unsigned(14 downto 0);
signal n7 : unsigned(14 downto 0);
signal n8 : unsigned(15 downto 0);
signal s9_1 : unsigned(14 downto 0);
component cf_ldpc_90 is
port (
i1 : in  unsigned(14 downto 0);
i2 : in  unsigned(14 downto 0);
i3 : in  unsigned(14 downto 0);
o1 : out unsigned(14 downto 0));
end component cf_ldpc_90;
begin
n1 <= i1(15 downto 15);
n2 <= i2(15 downto 15);
n3 <= i3(15 downto 15);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(14 downto 14) &
  i2(13 downto 13) &
  i2(12 downto 12) &
  i2(11 downto 11) &
  i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_90 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_88 is
port (
i1 : in  unsigned(16 downto 0);
i2 : in  unsigned(16 downto 0);
i3 : in  unsigned(16 downto 0);
o1 : out unsigned(16 downto 0));
end entity cf_ldpc_88;
architecture rtl of cf_ldpc_88 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(15 downto 0);
signal n6 : unsigned(15 downto 0);
signal n7 : unsigned(15 downto 0);
signal n8 : unsigned(16 downto 0);
signal s9_1 : unsigned(15 downto 0);
component cf_ldpc_89 is
port (
i1 : in  unsigned(15 downto 0);
i2 : in  unsigned(15 downto 0);
i3 : in  unsigned(15 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_ldpc_89;
begin
n1 <= i1(16 downto 16);
n2 <= i2(16 downto 16);
n3 <= i3(16 downto 16);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(15 downto 15) &
  i2(14 downto 14) &
  i2(13 downto 13) &
  i2(12 downto 12) &
  i2(11 downto 11) &
  i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_89 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_87 is
port (
i1 : in  unsigned(17 downto 0);
i2 : in  unsigned(17 downto 0);
i3 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end entity cf_ldpc_87;
architecture rtl of cf_ldpc_87 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(16 downto 0);
signal n6 : unsigned(16 downto 0);
signal n7 : unsigned(16 downto 0);
signal n8 : unsigned(17 downto 0);
signal s9_1 : unsigned(16 downto 0);
component cf_ldpc_88 is
port (
i1 : in  unsigned(16 downto 0);
i2 : in  unsigned(16 downto 0);
i3 : in  unsigned(16 downto 0);
o1 : out unsigned(16 downto 0));
end component cf_ldpc_88;
begin
n1 <= i1(17 downto 17);
n2 <= i2(17 downto 17);
n3 <= i3(17 downto 17);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(16 downto 16) &
  i2(15 downto 15) &
  i2(14 downto 14) &
  i2(13 downto 13) &
  i2(12 downto 12) &
  i2(11 downto 11) &
  i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_88 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_86 is
port (
i1 : in  unsigned(18 downto 0);
i2 : in  unsigned(18 downto 0);
i3 : in  unsigned(18 downto 0);
o1 : out unsigned(18 downto 0));
end entity cf_ldpc_86;
architecture rtl of cf_ldpc_86 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(17 downto 0);
signal n6 : unsigned(17 downto 0);
signal n7 : unsigned(17 downto 0);
signal n8 : unsigned(18 downto 0);
signal s9_1 : unsigned(17 downto 0);
component cf_ldpc_87 is
port (
i1 : in  unsigned(17 downto 0);
i2 : in  unsigned(17 downto 0);
i3 : in  unsigned(17 downto 0);
o1 : out unsigned(17 downto 0));
end component cf_ldpc_87;
begin
n1 <= i1(18 downto 18);
n2 <= i2(18 downto 18);
n3 <= i3(18 downto 18);
n4 <= n2 when n1 = "1" else n3;
n5 <= i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n6 <= i2(17 downto 17) &
  i2(16 downto 16) &
  i2(15 downto 15) &
  i2(14 downto 14) &
  i2(13 downto 13) &
  i2(12 downto 12) &
  i2(11 downto 11) &
  i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n7 <= i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_87 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_85 is
port (
i1 : in  unsigned(19 downto 0);
i2 : in  unsigned(19 downto 0);
i3 : in  unsigned(19 downto 0);
o1 : out unsigned(19 downto 0));
end entity cf_ldpc_85;
architecture rtl of cf_ldpc_85 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(18 downto 0);
signal n6 : unsigned(18 downto 0);
signal n7 : unsigned(18 downto 0);
signal n8 : unsigned(19 downto 0);
signal s9_1 : unsigned(18 downto 0);
component cf_ldpc_86 is
port (
i1 : in  unsigned(18 downto 0);
i2 : in  unsigned(18 downto 0);
i3 : in  unsigned(18 downto 0);
o1 : out unsigned(18 downto 0));
end component cf_ldpc_86;
begin
n1 <= i2(19 downto 19);
n2 <= i3(19 downto 19);
n3 <= i1(19 downto 19);
n4 <= n2 when n1 = "1" else n3;
n5 <= i2(18 downto 18) &
  i2(17 downto 17) &
  i2(16 downto 16) &
  i2(15 downto 15) &
  i2(14 downto 14) &
  i2(13 downto 13) &
  i2(12 downto 12) &
  i2(11 downto 11) &
  i2(10 downto 10) &
  i2(9 downto 9) &
  i2(8 downto 8) &
  i2(7 downto 7) &
  i2(6 downto 6) &
  i2(5 downto 5) &
  i2(4 downto 4) &
  i2(3 downto 3) &
  i2(2 downto 2) &
  i2(1 downto 1) &
  i2(0 downto 0);
n6 <= i3(18 downto 18) &
  i3(17 downto 17) &
  i3(16 downto 16) &
  i3(15 downto 15) &
  i3(14 downto 14) &
  i3(13 downto 13) &
  i3(12 downto 12) &
  i3(11 downto 11) &
  i3(10 downto 10) &
  i3(9 downto 9) &
  i3(8 downto 8) &
  i3(7 downto 7) &
  i3(6 downto 6) &
  i3(5 downto 5) &
  i3(4 downto 4) &
  i3(3 downto 3) &
  i3(2 downto 2) &
  i3(1 downto 1) &
  i3(0 downto 0);
n7 <= i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n8 <= n4 & s9_1;
s9 : cf_ldpc_86 port map (n5, n6, n7, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_84 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_ldpc_84;
architecture rtl of cf_ldpc_84 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
begin
n1 <= i1(15 downto 15) &
  i1(10 downto 10) &
  i1(5 downto 5);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_83 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(1 downto 0));
end entity cf_ldpc_83;
architecture rtl of cf_ldpc_83 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(1 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_ldpc_84 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_84;
begin
n1 <= i1(12 downto 12) &
  i1(8 downto 8) &
  i1(4 downto 4);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_84 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_82 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(2 downto 0));
end entity cf_ldpc_82;
architecture rtl of cf_ldpc_82 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(2 downto 0);
signal s10_1 : unsigned(1 downto 0);
component cf_ldpc_83 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(1 downto 0));
end component cf_ldpc_83;
begin
n1 <= i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_83 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_81 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(3 downto 0));
end entity cf_ldpc_81;
architecture rtl of cf_ldpc_81 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(3 downto 0);
signal s10_1 : unsigned(2 downto 0);
component cf_ldpc_82 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(2 downto 0));
end component cf_ldpc_82;
begin
n1 <= i1(17 downto 17) &
  i1(12 downto 12) &
  i1(7 downto 7);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_82 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_80 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(4 downto 0));
end entity cf_ldpc_80;
architecture rtl of cf_ldpc_80 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(4 downto 0);
signal s10_1 : unsigned(3 downto 0);
component cf_ldpc_81 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(3 downto 0));
end component cf_ldpc_81;
begin
n1 <= i1(16 downto 16) &
  i1(9 downto 9) &
  i1(5 downto 5);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_81 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_79 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(5 downto 0));
end entity cf_ldpc_79;
architecture rtl of cf_ldpc_79 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(5 downto 0);
signal s10_1 : unsigned(4 downto 0);
component cf_ldpc_80 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(4 downto 0));
end component cf_ldpc_80;
begin
n1 <= i1(3 downto 3) &
  i1(2 downto 2) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_80 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_78 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(6 downto 0));
end entity cf_ldpc_78;
architecture rtl of cf_ldpc_78 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(6 downto 0);
signal s10_1 : unsigned(5 downto 0);
component cf_ldpc_79 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(5 downto 0));
end component cf_ldpc_79;
begin
n1 <= i1(19 downto 19) &
  i1(14 downto 14) &
  i1(8 downto 8);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_79 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_77 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(7 downto 0));
end entity cf_ldpc_77;
architecture rtl of cf_ldpc_77 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(7 downto 0);
signal s10_1 : unsigned(6 downto 0);
component cf_ldpc_78 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(6 downto 0));
end component cf_ldpc_78;
begin
n1 <= i1(17 downto 17) &
  i1(13 downto 13) &
  i1(6 downto 6);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_78 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_76 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(8 downto 0));
end entity cf_ldpc_76;
architecture rtl of cf_ldpc_76 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(8 downto 0);
signal s10_1 : unsigned(7 downto 0);
component cf_ldpc_77 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(7 downto 0));
end component cf_ldpc_77;
begin
n1 <= i1(3 downto 3) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_77 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_75 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(9 downto 0));
end entity cf_ldpc_75;
architecture rtl of cf_ldpc_75 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(9 downto 0);
signal s10_1 : unsigned(8 downto 0);
component cf_ldpc_76 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_ldpc_76;
begin
n1 <= i1(16 downto 16) &
  i1(11 downto 11) &
  i1(6 downto 6);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_76 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_74 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(10 downto 0));
end entity cf_ldpc_74;
architecture rtl of cf_ldpc_74 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(10 downto 0);
signal s10_1 : unsigned(9 downto 0);
component cf_ldpc_75 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(9 downto 0));
end component cf_ldpc_75;
begin
n1 <= i1(18 downto 18) &
  i1(14 downto 14) &
  i1(10 downto 10);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_75 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_73 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(11 downto 0));
end entity cf_ldpc_73;
architecture rtl of cf_ldpc_73 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(11 downto 0);
signal s10_1 : unsigned(10 downto 0);
component cf_ldpc_74 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(10 downto 0));
end component cf_ldpc_74;
begin
n1 <= i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_74 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_72 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(12 downto 0));
end entity cf_ldpc_72;
architecture rtl of cf_ldpc_72 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(12 downto 0);
signal s10_1 : unsigned(11 downto 0);
component cf_ldpc_73 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(11 downto 0));
end component cf_ldpc_73;
begin
n1 <= i1(18 downto 18) &
  i1(13 downto 13) &
  i1(9 downto 9);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_73 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_71 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(13 downto 0));
end entity cf_ldpc_71;
architecture rtl of cf_ldpc_71 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(13 downto 0);
signal s10_1 : unsigned(12 downto 0);
component cf_ldpc_72 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(12 downto 0));
end component cf_ldpc_72;
begin
n1 <= i1(12 downto 12) &
  i1(8 downto 8) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_72 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_70 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(14 downto 0));
end entity cf_ldpc_70;
architecture rtl of cf_ldpc_70 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(14 downto 0);
signal s10_1 : unsigned(13 downto 0);
component cf_ldpc_71 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(13 downto 0));
end component cf_ldpc_71;
begin
n1 <= i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_71 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_69 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(15 downto 0));
end entity cf_ldpc_69;
architecture rtl of cf_ldpc_69 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(15 downto 0);
signal s10_1 : unsigned(14 downto 0);
component cf_ldpc_70 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(14 downto 0));
end component cf_ldpc_70;
begin
n1 <= i1(15 downto 15) &
  i1(10 downto 10) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_70 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_68 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(16 downto 0));
end entity cf_ldpc_68;
architecture rtl of cf_ldpc_68 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(16 downto 0);
signal s10_1 : unsigned(15 downto 0);
component cf_ldpc_69 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(15 downto 0));
end component cf_ldpc_69;
begin
n1 <= i1(16 downto 16) &
  i1(9 downto 9) &
  i1(1 downto 1);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_69 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_67 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(17 downto 0));
end entity cf_ldpc_67;
architecture rtl of cf_ldpc_67 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(17 downto 0);
signal s10_1 : unsigned(16 downto 0);
component cf_ldpc_68 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(16 downto 0));
end component cf_ldpc_68;
begin
n1 <= i1(7 downto 7) &
  i1(6 downto 6) &
  i1(4 downto 4);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_68 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_66 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(18 downto 0));
end entity cf_ldpc_66;
architecture rtl of cf_ldpc_66 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(18 downto 0);
signal s10_1 : unsigned(17 downto 0);
component cf_ldpc_67 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(17 downto 0));
end component cf_ldpc_67;
begin
n1 <= i1(16 downto 16) &
  i1(11 downto 11) &
  i1(3 downto 3);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_67 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_65 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(19 downto 0));
end entity cf_ldpc_65;
architecture rtl of cf_ldpc_65 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(19 downto 0);
signal s10_1 : unsigned(18 downto 0);
component cf_ldpc_66 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(18 downto 0));
end component cf_ldpc_66;
begin
n1 <= i1(17 downto 17) &
  i1(13 downto 13) &
  i1(2 downto 2);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_66 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_64 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(20 downto 0));
end entity cf_ldpc_64;
architecture rtl of cf_ldpc_64 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(20 downto 0);
signal s10_1 : unsigned(19 downto 0);
component cf_ldpc_65 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(19 downto 0));
end component cf_ldpc_65;
begin
n1 <= i1(7 downto 7) &
  i1(5 downto 5) &
  i1(4 downto 4);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_65 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_63 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(21 downto 0));
end entity cf_ldpc_63;
architecture rtl of cf_ldpc_63 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(21 downto 0);
signal s10_1 : unsigned(20 downto 0);
component cf_ldpc_64 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(20 downto 0));
end component cf_ldpc_64;
begin
n1 <= i1(17 downto 17) &
  i1(12 downto 12) &
  i1(1 downto 1);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_64 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_62 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(22 downto 0));
end entity cf_ldpc_62;
architecture rtl of cf_ldpc_62 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(22 downto 0);
signal s10_1 : unsigned(21 downto 0);
component cf_ldpc_63 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(21 downto 0));
end component cf_ldpc_63;
begin
n1 <= i1(19 downto 19) &
  i1(15 downto 15) &
  i1(11 downto 11);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_63 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_61 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(23 downto 0));
end entity cf_ldpc_61;
architecture rtl of cf_ldpc_61 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(23 downto 0);
signal s10_1 : unsigned(22 downto 0);
component cf_ldpc_62 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(22 downto 0));
end component cf_ldpc_62;
begin
n1 <= i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_62 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_60 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(24 downto 0));
end entity cf_ldpc_60;
architecture rtl of cf_ldpc_60 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(24 downto 0);
signal s10_1 : unsigned(23 downto 0);
component cf_ldpc_61 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(23 downto 0));
end component cf_ldpc_61;
begin
n1 <= i1(19 downto 19) &
  i1(14 downto 14) &
  i1(2 downto 2);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_61 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_59 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(25 downto 0));
end entity cf_ldpc_59;
architecture rtl of cf_ldpc_59 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(25 downto 0);
signal s10_1 : unsigned(24 downto 0);
component cf_ldpc_60 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(24 downto 0));
end component cf_ldpc_60;
begin
n1 <= i1(12 downto 12) &
  i1(4 downto 4) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_60 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_58 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(26 downto 0));
end entity cf_ldpc_58;
architecture rtl of cf_ldpc_58 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(26 downto 0);
signal s10_1 : unsigned(25 downto 0);
component cf_ldpc_59 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(25 downto 0));
end component cf_ldpc_59;
begin
n1 <= i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_59 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_57 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(27 downto 0));
end entity cf_ldpc_57;
architecture rtl of cf_ldpc_57 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(27 downto 0);
signal s10_1 : unsigned(26 downto 0);
component cf_ldpc_58 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(26 downto 0));
end component cf_ldpc_58;
begin
n1 <= i1(18 downto 18) &
  i1(13 downto 13) &
  i1(4 downto 4);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_58 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_56 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(28 downto 0));
end entity cf_ldpc_56;
architecture rtl of cf_ldpc_56 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(28 downto 0);
signal s10_1 : unsigned(27 downto 0);
component cf_ldpc_57 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(27 downto 0));
end component cf_ldpc_57;
begin
n1 <= i1(16 downto 16) &
  i1(5 downto 5) &
  i1(1 downto 1);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_57 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_55 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(29 downto 0));
end entity cf_ldpc_55;
architecture rtl of cf_ldpc_55 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(29 downto 0);
signal s10_1 : unsigned(28 downto 0);
component cf_ldpc_56 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(28 downto 0));
end component cf_ldpc_56;
begin
n1 <= i1(11 downto 11) &
  i1(10 downto 10) &
  i1(8 downto 8);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_56 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_54 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(30 downto 0));
end entity cf_ldpc_54;
architecture rtl of cf_ldpc_54 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(30 downto 0);
signal s10_1 : unsigned(29 downto 0);
component cf_ldpc_55 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(29 downto 0));
end component cf_ldpc_55;
begin
n1 <= i1(15 downto 15) &
  i1(5 downto 5) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_55 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_53 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(31 downto 0));
end entity cf_ldpc_53;
architecture rtl of cf_ldpc_53 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(31 downto 0);
signal s10_1 : unsigned(30 downto 0);
component cf_ldpc_54 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(30 downto 0));
end component cf_ldpc_54;
begin
n1 <= i1(18 downto 18) &
  i1(14 downto 14) &
  i1(3 downto 3);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_54 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_52 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(32 downto 0));
end entity cf_ldpc_52;
architecture rtl of cf_ldpc_52 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(32 downto 0);
signal s10_1 : unsigned(31 downto 0);
component cf_ldpc_53 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(31 downto 0));
end component cf_ldpc_53;
begin
n1 <= i1(11 downto 11) &
  i1(9 downto 9) &
  i1(8 downto 8);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_53 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_51 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(33 downto 0));
end entity cf_ldpc_51;
architecture rtl of cf_ldpc_51 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(33 downto 0);
signal s10_1 : unsigned(32 downto 0);
component cf_ldpc_52 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(32 downto 0));
end component cf_ldpc_52;
begin
n1 <= i1(16 downto 16) &
  i1(6 downto 6) &
  i1(3 downto 3);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_52 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_50 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(34 downto 0));
end entity cf_ldpc_50;
architecture rtl of cf_ldpc_50 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(34 downto 0);
signal s10_1 : unsigned(33 downto 0);
component cf_ldpc_51 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(33 downto 0));
end component cf_ldpc_51;
begin
n1 <= i1(19 downto 19) &
  i1(15 downto 15) &
  i1(7 downto 7);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_51 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_49 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(35 downto 0));
end entity cf_ldpc_49;
architecture rtl of cf_ldpc_49 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(35 downto 0);
signal s10_1 : unsigned(34 downto 0);
component cf_ldpc_50 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(34 downto 0));
end component cf_ldpc_50;
begin
n1 <= i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_50 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_48 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(36 downto 0));
end entity cf_ldpc_48;
architecture rtl of cf_ldpc_48 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(36 downto 0);
signal s10_1 : unsigned(35 downto 0);
component cf_ldpc_49 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(35 downto 0));
end component cf_ldpc_49;
begin
n1 <= i1(17 downto 17) &
  i1(7 downto 7) &
  i1(1 downto 1);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_49 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_47 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(37 downto 0));
end entity cf_ldpc_47;
architecture rtl of cf_ldpc_47 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(37 downto 0);
signal s10_1 : unsigned(36 downto 0);
component cf_ldpc_48 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(36 downto 0));
end component cf_ldpc_48;
begin
n1 <= i1(8 downto 8) &
  i1(4 downto 4) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_48 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_46 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(38 downto 0));
end entity cf_ldpc_46;
architecture rtl of cf_ldpc_46 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(38 downto 0);
signal s10_1 : unsigned(37 downto 0);
component cf_ldpc_47 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(37 downto 0));
end component cf_ldpc_47;
begin
n1 <= i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_47 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_45 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(39 downto 0));
end entity cf_ldpc_45;
architecture rtl of cf_ldpc_45 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(39 downto 0);
signal s10_1 : unsigned(38 downto 0);
component cf_ldpc_46 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(38 downto 0));
end component cf_ldpc_46;
begin
n1 <= i1(18 downto 18) &
  i1(9 downto 9) &
  i1(4 downto 4);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_46 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_44 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(40 downto 0));
end entity cf_ldpc_44;
architecture rtl of cf_ldpc_44 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(40 downto 0);
signal s10_1 : unsigned(39 downto 0);
component cf_ldpc_45 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(39 downto 0));
end component cf_ldpc_45;
begin
n1 <= i1(17 downto 17) &
  i1(6 downto 6) &
  i1(2 downto 2);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_45 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_43 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(41 downto 0));
end entity cf_ldpc_43;
architecture rtl of cf_ldpc_43 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(41 downto 0);
signal s10_1 : unsigned(40 downto 0);
component cf_ldpc_44 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(40 downto 0));
end component cf_ldpc_44;
begin
n1 <= i1(15 downto 15) &
  i1(14 downto 14) &
  i1(12 downto 12);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_44 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_42 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(42 downto 0));
end entity cf_ldpc_42;
architecture rtl of cf_ldpc_42 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(42 downto 0);
signal s10_1 : unsigned(41 downto 0);
component cf_ldpc_43 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(41 downto 0));
end component cf_ldpc_43;
begin
n1 <= i1(19 downto 19) &
  i1(8 downto 8) &
  i1(2 downto 2);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_43 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_41 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(43 downto 0));
end entity cf_ldpc_41;
architecture rtl of cf_ldpc_41 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(43 downto 0);
signal s10_1 : unsigned(42 downto 0);
component cf_ldpc_42 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(42 downto 0));
end component cf_ldpc_42;
begin
n1 <= i1(18 downto 18) &
  i1(10 downto 10) &
  i1(3 downto 3);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_42 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_40 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(44 downto 0));
end entity cf_ldpc_40;
architecture rtl of cf_ldpc_40 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(44 downto 0);
signal s10_1 : unsigned(43 downto 0);
component cf_ldpc_41 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(43 downto 0));
end component cf_ldpc_41;
begin
n1 <= i1(15 downto 15) &
  i1(13 downto 13) &
  i1(12 downto 12);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_41 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_39 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(45 downto 0));
end entity cf_ldpc_39;
architecture rtl of cf_ldpc_39 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(45 downto 0);
signal s10_1 : unsigned(44 downto 0);
component cf_ldpc_40 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(44 downto 0));
end component cf_ldpc_40;
begin
n1 <= i1(10 downto 10) &
  i1(5 downto 5) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_40 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_38 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(46 downto 0));
end entity cf_ldpc_38;
architecture rtl of cf_ldpc_38 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(46 downto 0);
signal s10_1 : unsigned(45 downto 0);
component cf_ldpc_39 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(45 downto 0));
end component cf_ldpc_39;
begin
n1 <= i1(19 downto 19) &
  i1(11 downto 11) &
  i1(7 downto 7);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_39 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_37 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(47 downto 0));
end entity cf_ldpc_37;
architecture rtl of cf_ldpc_37 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(47 downto 0);
signal s10_1 : unsigned(46 downto 0);
component cf_ldpc_38 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(46 downto 0));
end component cf_ldpc_38;
begin
n1 <= i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_38 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_36 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(48 downto 0));
end entity cf_ldpc_36;
architecture rtl of cf_ldpc_36 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(48 downto 0);
signal s10_1 : unsigned(47 downto 0);
component cf_ldpc_37 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(47 downto 0));
end component cf_ldpc_37;
begin
n1 <= i1(11 downto 11) &
  i1(6 downto 6) &
  i1(3 downto 3);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_37 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_35 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(49 downto 0));
end entity cf_ldpc_35;
architecture rtl of cf_ldpc_35 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(49 downto 0);
signal s10_1 : unsigned(48 downto 0);
component cf_ldpc_36 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(48 downto 0));
end component cf_ldpc_36;
begin
n1 <= i1(9 downto 9) &
  i1(5 downto 5) &
  i1(1 downto 1);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_36 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_34 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(50 downto 0));
end entity cf_ldpc_34;
architecture rtl of cf_ldpc_34 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(50 downto 0);
signal s10_1 : unsigned(49 downto 0);
component cf_ldpc_35 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(49 downto 0));
end component cf_ldpc_35;
begin
n1 <= i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_35 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_33 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(51 downto 0));
end entity cf_ldpc_33;
architecture rtl of cf_ldpc_33 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(51 downto 0);
signal s10_1 : unsigned(50 downto 0);
component cf_ldpc_34 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(50 downto 0));
end component cf_ldpc_34;
begin
n1 <= i1(12 downto 12) &
  i1(7 downto 7) &
  i1(1 downto 1);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_34 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_32 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(52 downto 0));
end entity cf_ldpc_32;
architecture rtl of cf_ldpc_32 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(52 downto 0);
signal s10_1 : unsigned(51 downto 0);
component cf_ldpc_33 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(51 downto 0));
end component cf_ldpc_33;
begin
n1 <= i1(13 downto 13) &
  i1(6 downto 6) &
  i1(2 downto 2);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_33 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_31 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(53 downto 0));
end entity cf_ldpc_31;
architecture rtl of cf_ldpc_31 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(53 downto 0);
signal s10_1 : unsigned(52 downto 0);
component cf_ldpc_32 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(52 downto 0));
end component cf_ldpc_32;
begin
n1 <= i1(19 downto 19) &
  i1(18 downto 18) &
  i1(16 downto 16);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_32 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_30 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(54 downto 0));
end entity cf_ldpc_30;
architecture rtl of cf_ldpc_30 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(54 downto 0);
signal s10_1 : unsigned(53 downto 0);
component cf_ldpc_31 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(53 downto 0));
end component cf_ldpc_31;
begin
n1 <= i1(13 downto 13) &
  i1(9 downto 9) &
  i1(4 downto 4);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_31 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_29 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(55 downto 0));
end entity cf_ldpc_29;
architecture rtl of cf_ldpc_29 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(55 downto 0);
signal s10_1 : unsigned(54 downto 0);
component cf_ldpc_30 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(54 downto 0));
end component cf_ldpc_30;
begin
n1 <= i1(14 downto 14) &
  i1(10 downto 10) &
  i1(3 downto 3);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_30 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_28 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(56 downto 0));
end entity cf_ldpc_28;
architecture rtl of cf_ldpc_28 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(56 downto 0);
signal s10_1 : unsigned(55 downto 0);
component cf_ldpc_29 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(55 downto 0));
end component cf_ldpc_29;
begin
n1 <= i1(19 downto 19) &
  i1(17 downto 17) &
  i1(16 downto 16);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_29 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_27 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(57 downto 0));
end entity cf_ldpc_27;
architecture rtl of cf_ldpc_27 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(57 downto 0);
signal s10_1 : unsigned(56 downto 0);
component cf_ldpc_28 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(56 downto 0));
end component cf_ldpc_28;
begin
n1 <= i1(14 downto 14) &
  i1(8 downto 8) &
  i1(2 downto 2);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_28 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_26 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(58 downto 0));
end entity cf_ldpc_26;
architecture rtl of cf_ldpc_26 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(58 downto 0);
signal s10_1 : unsigned(57 downto 0);
component cf_ldpc_27 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(57 downto 0));
end component cf_ldpc_27;
begin
n1 <= i1(15 downto 15) &
  i1(11 downto 11) &
  i1(7 downto 7);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_27 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_25 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(59 downto 0));
end entity cf_ldpc_25;
architecture rtl of cf_ldpc_25 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(1 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(59 downto 0);
signal s10_1 : unsigned(58 downto 0);
component cf_ldpc_26 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(58 downto 0));
end component cf_ldpc_26;
begin
n1 <= i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16);
n2 <= n1(2 downto 2);
n3 <= n1(1 downto 1) &
  n1(0 downto 0);
n4 <= n3(1 downto 1);
n5 <= n3(0 downto 0);
n6 <= n5(0 downto 0);
n7 <= n2 xor n4;
n8 <= n7 xor n6;
n9 <= n8 & s10_1;
s10 : cf_ldpc_26 port map (i1, s10_1);
o1 <= n9;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_24 is
port (
i1 : in  unsigned(4 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0));
end entity cf_ldpc_24;
architecture rtl of cf_ldpc_24 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(3 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(2 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(1 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
begin
n1 <= i1(4 downto 4);
n2 <= i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n3 <= n2(3 downto 3);
n4 <= n2(2 downto 2) &
  n2(1 downto 1) &
  n2(0 downto 0);
n5 <= n4(2 downto 2);
n6 <= n4(1 downto 1) &
  n4(0 downto 0);
n7 <= n6(1 downto 1);
n8 <= n6(0 downto 0);
n9 <= n8(0 downto 0);
o5 <= n9;
o4 <= n7;
o3 <= n5;
o2 <= n3;
o1 <= n1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_23 is
port (
i1 : in  unsigned(8 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0);
o9 : out unsigned(0 downto 0));
end entity cf_ldpc_23;
architecture rtl of cf_ldpc_23 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(7 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(6 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(5 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(4 downto 0);
signal s9_1 : unsigned(0 downto 0);
signal s9_2 : unsigned(0 downto 0);
signal s9_3 : unsigned(0 downto 0);
signal s9_4 : unsigned(0 downto 0);
signal s9_5 : unsigned(0 downto 0);
component cf_ldpc_24 is
port (
i1 : in  unsigned(4 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0));
end component cf_ldpc_24;
begin
n1 <= i1(8 downto 8);
n2 <= i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n3 <= n2(7 downto 7);
n4 <= n2(6 downto 6) &
  n2(5 downto 5) &
  n2(4 downto 4) &
  n2(3 downto 3) &
  n2(2 downto 2) &
  n2(1 downto 1) &
  n2(0 downto 0);
n5 <= n4(6 downto 6);
n6 <= n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
n7 <= n6(5 downto 5);
n8 <= n6(4 downto 4) &
  n6(3 downto 3) &
  n6(2 downto 2) &
  n6(1 downto 1) &
  n6(0 downto 0);
s9 : cf_ldpc_24 port map (n8, s9_1, s9_2, s9_3, s9_4, s9_5);
o9 <= s9_5;
o8 <= s9_4;
o7 <= s9_3;
o6 <= s9_2;
o5 <= s9_1;
o4 <= n7;
o3 <= n5;
o2 <= n3;
o1 <= n1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_22 is
port (
i1 : in  unsigned(12 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0);
o9 : out unsigned(0 downto 0);
o10 : out unsigned(0 downto 0);
o11 : out unsigned(0 downto 0);
o12 : out unsigned(0 downto 0);
o13 : out unsigned(0 downto 0));
end entity cf_ldpc_22;
architecture rtl of cf_ldpc_22 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(11 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(10 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(9 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(8 downto 0);
signal s9_1 : unsigned(0 downto 0);
signal s9_2 : unsigned(0 downto 0);
signal s9_3 : unsigned(0 downto 0);
signal s9_4 : unsigned(0 downto 0);
signal s9_5 : unsigned(0 downto 0);
signal s9_6 : unsigned(0 downto 0);
signal s9_7 : unsigned(0 downto 0);
signal s9_8 : unsigned(0 downto 0);
signal s9_9 : unsigned(0 downto 0);
component cf_ldpc_23 is
port (
i1 : in  unsigned(8 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0);
o9 : out unsigned(0 downto 0));
end component cf_ldpc_23;
begin
n1 <= i1(12 downto 12);
n2 <= i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n3 <= n2(11 downto 11);
n4 <= n2(10 downto 10) &
  n2(9 downto 9) &
  n2(8 downto 8) &
  n2(7 downto 7) &
  n2(6 downto 6) &
  n2(5 downto 5) &
  n2(4 downto 4) &
  n2(3 downto 3) &
  n2(2 downto 2) &
  n2(1 downto 1) &
  n2(0 downto 0);
n5 <= n4(10 downto 10);
n6 <= n4(9 downto 9) &
  n4(8 downto 8) &
  n4(7 downto 7) &
  n4(6 downto 6) &
  n4(5 downto 5) &
  n4(4 downto 4) &
  n4(3 downto 3) &
  n4(2 downto 2) &
  n4(1 downto 1) &
  n4(0 downto 0);
n7 <= n6(9 downto 9);
n8 <= n6(8 downto 8) &
  n6(7 downto 7) &
  n6(6 downto 6) &
  n6(5 downto 5) &
  n6(4 downto 4) &
  n6(3 downto 3) &
  n6(2 downto 2) &
  n6(1 downto 1) &
  n6(0 downto 0);
s9 : cf_ldpc_23 port map (n8, s9_1, s9_2, s9_3, s9_4, s9_5, s9_6, s9_7, s9_8, s9_9);
o13 <= s9_9;
o12 <= s9_8;
o11 <= s9_7;
o10 <= s9_6;
o9 <= s9_5;
o8 <= s9_4;
o7 <= s9_3;
o6 <= s9_2;
o5 <= s9_1;
o4 <= n7;
o3 <= n5;
o2 <= n3;
o1 <= n1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_21 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
i10 : in  unsigned(0 downto 0);
i11 : in  unsigned(0 downto 0);
i12 : in  unsigned(0 downto 0);
i13 : in  unsigned(0 downto 0);
i14 : in  unsigned(0 downto 0);
i15 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_ldpc_21;
architecture rtl of cf_ldpc_21 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
signal n11 : unsigned(0 downto 0);
signal n12 : unsigned(0 downto 0);
signal n13 : unsigned(0 downto 0);
signal n14 : unsigned(0 downto 0);
begin
n1 <= i1 or i2;
n2 <= i3 or i4;
n3 <= i5 or i6;
n4 <= i7 or i8;
n5 <= i9 or i10;
n6 <= i11 or i12;
n7 <= i13 or i14;
n8 <= n1 or n2;
n9 <= n3 or n4;
n10 <= n5 or n6;
n11 <= n7 or i15;
n12 <= n8 or n9;
n13 <= n10 or n11;
n14 <= n12 or n13;
o1 <= n14;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_20 is
port (
i1 : in  unsigned(3 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_ldpc_20;
architecture rtl of cf_ldpc_20 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(2 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(1 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(0 downto 0);
begin
n1 <= i1(3 downto 3);
n2 <= i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n3 <= n2(2 downto 2);
n4 <= n2(1 downto 1) &
  n2(0 downto 0);
n5 <= n4(1 downto 1);
n6 <= n4(0 downto 0);
n7 <= n6(0 downto 0);
n8 <= n1 xor n3;
n9 <= n5 xor n7;
n10 <= n8 xor n9;
o1 <= n10;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_19 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(2 downto 0));
end entity cf_ldpc_19;
architecture rtl of cf_ldpc_19 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(3 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(1 downto 0);
signal n5 : unsigned(2 downto 0);
signal s6_1 : unsigned(0 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_ldpc_20 is
port (
i1 : in  unsigned(3 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_20;
begin
n1 <= i1(17 downto 17) &
  i1(12 downto 12) &
  i1(7 downto 7) &
  i1(1 downto 1);
n2 <= i1(16 downto 16) &
  i1(11 downto 11) &
  i1(6 downto 6) &
  i1(3 downto 3);
n3 <= i1(15 downto 15) &
  i1(10 downto 10) &
  i1(5 downto 5) &
  i1(0 downto 0);
n4 <= s7_1 & s6_1;
n5 <= s8_1 & n4;
s6 : cf_ldpc_20 port map (n3, s6_1);
s7 : cf_ldpc_20 port map (n2, s7_1);
s8 : cf_ldpc_20 port map (n1, s8_1);
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_18 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(5 downto 0));
end entity cf_ldpc_18;
architecture rtl of cf_ldpc_18 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(3 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(3 downto 0);
signal n5 : unsigned(4 downto 0);
signal n6 : unsigned(5 downto 0);
signal s7_1 : unsigned(2 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s9_1 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_ldpc_19 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(2 downto 0));
end component cf_ldpc_19;
component cf_ldpc_20 is
port (
i1 : in  unsigned(3 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_20;
begin
n1 <= i1(12 downto 12) &
  i1(8 downto 8) &
  i1(4 downto 4) &
  i1(0 downto 0);
n2 <= i1(19 downto 19) &
  i1(14 downto 14) &
  i1(8 downto 8) &
  i1(2 downto 2);
n3 <= i1(18 downto 18) &
  i1(13 downto 13) &
  i1(9 downto 9) &
  i1(4 downto 4);
n4 <= s8_1 & s7_1;
n5 <= s9_1 & n4;
n6 <= s10_1 & n5;
s7 : cf_ldpc_19 port map (i1, s7_1);
s8 : cf_ldpc_20 port map (n3, s8_1);
s9 : cf_ldpc_20 port map (n2, s9_1);
s10 : cf_ldpc_20 port map (n1, s10_1);
o1 <= n6;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_17 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(8 downto 0));
end entity cf_ldpc_17;
architecture rtl of cf_ldpc_17 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(3 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(6 downto 0);
signal n5 : unsigned(7 downto 0);
signal n6 : unsigned(8 downto 0);
signal s7_1 : unsigned(5 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s9_1 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_ldpc_18 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(5 downto 0));
end component cf_ldpc_18;
component cf_ldpc_20 is
port (
i1 : in  unsigned(3 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_20;
begin
n1 <= i1(18 downto 18) &
  i1(14 downto 14) &
  i1(10 downto 10) &
  i1(3 downto 3);
n2 <= i1(17 downto 17) &
  i1(13 downto 13) &
  i1(6 downto 6) &
  i1(2 downto 2);
n3 <= i1(16 downto 16) &
  i1(9 downto 9) &
  i1(5 downto 5) &
  i1(1 downto 1);
n4 <= s8_1 & s7_1;
n5 <= s9_1 & n4;
n6 <= s10_1 & n5;
s7 : cf_ldpc_18 port map (i1, s7_1);
s8 : cf_ldpc_20 port map (n3, s8_1);
s9 : cf_ldpc_20 port map (n2, s9_1);
s10 : cf_ldpc_20 port map (n1, s10_1);
o1 <= n6;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_16 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(11 downto 0));
end entity cf_ldpc_16;
architecture rtl of cf_ldpc_16 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(3 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(9 downto 0);
signal n5 : unsigned(10 downto 0);
signal n6 : unsigned(11 downto 0);
signal s7_1 : unsigned(8 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s9_1 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_ldpc_17 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(8 downto 0));
end component cf_ldpc_17;
component cf_ldpc_20 is
port (
i1 : in  unsigned(3 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_20;
begin
n1 <= i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4);
n2 <= i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n3 <= i1(19 downto 19) &
  i1(15 downto 15) &
  i1(11 downto 11) &
  i1(7 downto 7);
n4 <= s8_1 & s7_1;
n5 <= s9_1 & n4;
n6 <= s10_1 & n5;
s7 : cf_ldpc_17 port map (i1, s7_1);
s8 : cf_ldpc_20 port map (n3, s8_1);
s9 : cf_ldpc_20 port map (n2, s9_1);
s10 : cf_ldpc_20 port map (n1, s10_1);
o1 <= n6;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_15 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(14 downto 0));
end entity cf_ldpc_15;
architecture rtl of cf_ldpc_15 is
signal n1 : unsigned(3 downto 0);
signal n2 : unsigned(3 downto 0);
signal n3 : unsigned(3 downto 0);
signal n4 : unsigned(12 downto 0);
signal n5 : unsigned(13 downto 0);
signal n6 : unsigned(14 downto 0);
signal s7_1 : unsigned(11 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s9_1 : unsigned(0 downto 0);
signal s10_1 : unsigned(0 downto 0);
component cf_ldpc_16 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(11 downto 0));
end component cf_ldpc_16;
component cf_ldpc_20 is
port (
i1 : in  unsigned(3 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_20;
begin
n1 <= i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16);
n2 <= i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12);
n3 <= i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8);
n4 <= s8_1 & s7_1;
n5 <= s9_1 & n4;
n6 <= s10_1 & n5;
s7 : cf_ldpc_16 port map (i1, s7_1);
s8 : cf_ldpc_20 port map (n3, s8_1);
s9 : cf_ldpc_20 port map (n2, s9_1);
s10 : cf_ldpc_20 port map (n1, s10_1);
o1 <= n6;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_14 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_ldpc_14;
architecture rtl of cf_ldpc_14 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(13 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(12 downto 0);
signal n5 : unsigned(0 downto 0);
signal s6_1 : unsigned(0 downto 0);
signal s6_2 : unsigned(0 downto 0);
signal s6_3 : unsigned(0 downto 0);
signal s6_4 : unsigned(0 downto 0);
signal s6_5 : unsigned(0 downto 0);
signal s6_6 : unsigned(0 downto 0);
signal s6_7 : unsigned(0 downto 0);
signal s6_8 : unsigned(0 downto 0);
signal s6_9 : unsigned(0 downto 0);
signal s6_10 : unsigned(0 downto 0);
signal s6_11 : unsigned(0 downto 0);
signal s6_12 : unsigned(0 downto 0);
signal s6_13 : unsigned(0 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s8_1 : unsigned(14 downto 0);
component cf_ldpc_22 is
port (
i1 : in  unsigned(12 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(0 downto 0);
o3 : out unsigned(0 downto 0);
o4 : out unsigned(0 downto 0);
o5 : out unsigned(0 downto 0);
o6 : out unsigned(0 downto 0);
o7 : out unsigned(0 downto 0);
o8 : out unsigned(0 downto 0);
o9 : out unsigned(0 downto 0);
o10 : out unsigned(0 downto 0);
o11 : out unsigned(0 downto 0);
o12 : out unsigned(0 downto 0);
o13 : out unsigned(0 downto 0));
end component cf_ldpc_22;
component cf_ldpc_21 is
port (
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(0 downto 0);
i3 : in  unsigned(0 downto 0);
i4 : in  unsigned(0 downto 0);
i5 : in  unsigned(0 downto 0);
i6 : in  unsigned(0 downto 0);
i7 : in  unsigned(0 downto 0);
i8 : in  unsigned(0 downto 0);
i9 : in  unsigned(0 downto 0);
i10 : in  unsigned(0 downto 0);
i11 : in  unsigned(0 downto 0);
i12 : in  unsigned(0 downto 0);
i13 : in  unsigned(0 downto 0);
i14 : in  unsigned(0 downto 0);
i15 : in  unsigned(0 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_21;
component cf_ldpc_15 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(14 downto 0));
end component cf_ldpc_15;
begin
n1 <= s8_1(14 downto 14);
n2 <= s8_1(13 downto 13) &
  s8_1(12 downto 12) &
  s8_1(11 downto 11) &
  s8_1(10 downto 10) &
  s8_1(9 downto 9) &
  s8_1(8 downto 8) &
  s8_1(7 downto 7) &
  s8_1(6 downto 6) &
  s8_1(5 downto 5) &
  s8_1(4 downto 4) &
  s8_1(3 downto 3) &
  s8_1(2 downto 2) &
  s8_1(1 downto 1) &
  s8_1(0 downto 0);
n3 <= n2(13 downto 13);
n4 <= n2(12 downto 12) &
  n2(11 downto 11) &
  n2(10 downto 10) &
  n2(9 downto 9) &
  n2(8 downto 8) &
  n2(7 downto 7) &
  n2(6 downto 6) &
  n2(5 downto 5) &
  n2(4 downto 4) &
  n2(3 downto 3) &
  n2(2 downto 2) &
  n2(1 downto 1) &
  n2(0 downto 0);
n5 <= not s7_1;
s6 : cf_ldpc_22 port map (n4, s6_1, s6_2, s6_3, s6_4, s6_5, s6_6, s6_7, s6_8, s6_9, s6_10, s6_11, s6_12, s6_13);
s7 : cf_ldpc_21 port map (n1, n3, s6_1, s6_2, s6_3, s6_4, s6_5, s6_6, s6_7, s6_8, s6_9, s6_10, s6_11, s6_12, s6_13, s7_1);
s8 : cf_ldpc_15 port map (i1, s8_1);
o1 <= n5;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_13 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_ldpc_13;
architecture rtl of cf_ldpc_13 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
begin
n1 <= i1(2 downto 2);
n2 <= i1(1 downto 1) &
  i1(0 downto 0);
n3 <= n2(1 downto 1);
n4 <= n2(0 downto 0);
n5 <= n4(0 downto 0);
n6 <= n1 or n3;
n7 <= n6 or n5;
n8 <= not n7;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end entity cf_ldpc_12;
architecture rtl of cf_ldpc_12 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(1 downto 0);
signal n3 : unsigned(0 downto 0);
signal n4 : unsigned(0 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(0 downto 0);
signal n7 : unsigned(0 downto 0);
signal n8 : unsigned(0 downto 0);
signal s9_1 : unsigned(0 downto 0);
component cf_ldpc_13 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_13;
begin
n1 <= i1(2 downto 2);
n2 <= i1(1 downto 1) &
  i1(0 downto 0);
n3 <= n2(1 downto 1);
n4 <= n2(0 downto 0);
n5 <= n4(0 downto 0);
n6 <= n1 and n3;
n7 <= n6 and n5;
n8 <= n7 or s9_1;
s9 : cf_ldpc_13 port map (i1, s9_1);
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_11 is
port (
i1 : in  unsigned(5 downto 0);
o1 : out unsigned(1 downto 0);
o2 : out unsigned(1 downto 0));
end entity cf_ldpc_11;
architecture rtl of cf_ldpc_11 is
signal n1 : unsigned(2 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(1 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(1 downto 0);
signal s7_1 : unsigned(0 downto 0);
signal s8_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
begin
n1 <= i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(2 downto 2);
n3 <= i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3);
n4 <= s8_1 & s7_1;
n5 <= i1(5 downto 5);
n6 <= n5 & n2;
s7 : cf_ldpc_12 port map (n1, s7_1);
s8 : cf_ldpc_12 port map (n3, s8_1);
o2 <= n6;
o1 <= n4;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_10 is
port (
i1 : in  unsigned(11 downto 0);
o1 : out unsigned(3 downto 0);
o2 : out unsigned(3 downto 0));
end entity cf_ldpc_10;
architecture rtl of cf_ldpc_10 is
signal n1 : unsigned(8 downto 0);
signal n2 : unsigned(5 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(2 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(2 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(3 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(3 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(1 downto 0);
signal s12_2 : unsigned(1 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_11 is
port (
i1 : in  unsigned(5 downto 0);
o1 : out unsigned(1 downto 0);
o2 : out unsigned(1 downto 0));
end component cf_ldpc_11;
begin
n1 <= i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6);
n4 <= s11_1 & s12_1;
n5 <= n1(8 downto 8);
n6 <= n5 & s12_2;
n7 <= i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9);
n8 <= s13_1 & n4;
n9 <= i1(11 downto 11);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_11 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_9 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(5 downto 0);
o2 : out unsigned(5 downto 0));
end entity cf_ldpc_9;
architecture rtl of cf_ldpc_9 is
signal n1 : unsigned(14 downto 0);
signal n2 : unsigned(11 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(4 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(4 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(5 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(5 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(3 downto 0);
signal s12_2 : unsigned(3 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_10 is
port (
i1 : in  unsigned(11 downto 0);
o1 : out unsigned(3 downto 0);
o2 : out unsigned(3 downto 0));
end component cf_ldpc_10;
begin
n1 <= i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12);
n4 <= s11_1 & s12_1;
n5 <= n1(14 downto 14);
n6 <= n5 & s12_2;
n7 <= i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15);
n8 <= s13_1 & n4;
n9 <= i1(17 downto 17);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_10 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_8 is
port (
i1 : in  unsigned(23 downto 0);
o1 : out unsigned(7 downto 0);
o2 : out unsigned(7 downto 0));
end entity cf_ldpc_8;
architecture rtl of cf_ldpc_8 is
signal n1 : unsigned(20 downto 0);
signal n2 : unsigned(17 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(6 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(6 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(7 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(7 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(5 downto 0);
signal s12_2 : unsigned(5 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_9 is
port (
i1 : in  unsigned(17 downto 0);
o1 : out unsigned(5 downto 0);
o2 : out unsigned(5 downto 0));
end component cf_ldpc_9;
begin
n1 <= i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18);
n4 <= s11_1 & s12_1;
n5 <= n1(20 downto 20);
n6 <= n5 & s12_2;
n7 <= i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21);
n8 <= s13_1 & n4;
n9 <= i1(23 downto 23);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_9 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_7 is
port (
i1 : in  unsigned(29 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(9 downto 0));
end entity cf_ldpc_7;
architecture rtl of cf_ldpc_7 is
signal n1 : unsigned(26 downto 0);
signal n2 : unsigned(23 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(8 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(8 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(9 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(9 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(7 downto 0);
signal s12_2 : unsigned(7 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_8 is
port (
i1 : in  unsigned(23 downto 0);
o1 : out unsigned(7 downto 0);
o2 : out unsigned(7 downto 0));
end component cf_ldpc_8;
begin
n1 <= i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24);
n4 <= s11_1 & s12_1;
n5 <= n1(26 downto 26);
n6 <= n5 & s12_2;
n7 <= i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27);
n8 <= s13_1 & n4;
n9 <= i1(29 downto 29);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_8 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_6 is
port (
i1 : in  unsigned(35 downto 0);
o1 : out unsigned(11 downto 0);
o2 : out unsigned(11 downto 0));
end entity cf_ldpc_6;
architecture rtl of cf_ldpc_6 is
signal n1 : unsigned(32 downto 0);
signal n2 : unsigned(29 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(10 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(10 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(11 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(11 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(9 downto 0);
signal s12_2 : unsigned(9 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_7 is
port (
i1 : in  unsigned(29 downto 0);
o1 : out unsigned(9 downto 0);
o2 : out unsigned(9 downto 0));
end component cf_ldpc_7;
begin
n1 <= i1(32 downto 32) &
  i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30);
n4 <= s11_1 & s12_1;
n5 <= n1(32 downto 32);
n6 <= n5 & s12_2;
n7 <= i1(35 downto 35) &
  i1(34 downto 34) &
  i1(33 downto 33);
n8 <= s13_1 & n4;
n9 <= i1(35 downto 35);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_7 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_5 is
port (
i1 : in  unsigned(41 downto 0);
o1 : out unsigned(13 downto 0);
o2 : out unsigned(13 downto 0));
end entity cf_ldpc_5;
architecture rtl of cf_ldpc_5 is
signal n1 : unsigned(38 downto 0);
signal n2 : unsigned(35 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(12 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(12 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(13 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(13 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(11 downto 0);
signal s12_2 : unsigned(11 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_6 is
port (
i1 : in  unsigned(35 downto 0);
o1 : out unsigned(11 downto 0);
o2 : out unsigned(11 downto 0));
end component cf_ldpc_6;
begin
n1 <= i1(38 downto 38) &
  i1(37 downto 37) &
  i1(36 downto 36) &
  i1(35 downto 35) &
  i1(34 downto 34) &
  i1(33 downto 33) &
  i1(32 downto 32) &
  i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(38 downto 38) &
  n1(37 downto 37) &
  n1(36 downto 36);
n4 <= s11_1 & s12_1;
n5 <= n1(38 downto 38);
n6 <= n5 & s12_2;
n7 <= i1(41 downto 41) &
  i1(40 downto 40) &
  i1(39 downto 39);
n8 <= s13_1 & n4;
n9 <= i1(41 downto 41);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_6 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_4 is
port (
i1 : in  unsigned(47 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end entity cf_ldpc_4;
architecture rtl of cf_ldpc_4 is
signal n1 : unsigned(44 downto 0);
signal n2 : unsigned(41 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(14 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(14 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(15 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(15 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(13 downto 0);
signal s12_2 : unsigned(13 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_5 is
port (
i1 : in  unsigned(41 downto 0);
o1 : out unsigned(13 downto 0);
o2 : out unsigned(13 downto 0));
end component cf_ldpc_5;
begin
n1 <= i1(44 downto 44) &
  i1(43 downto 43) &
  i1(42 downto 42) &
  i1(41 downto 41) &
  i1(40 downto 40) &
  i1(39 downto 39) &
  i1(38 downto 38) &
  i1(37 downto 37) &
  i1(36 downto 36) &
  i1(35 downto 35) &
  i1(34 downto 34) &
  i1(33 downto 33) &
  i1(32 downto 32) &
  i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(41 downto 41) &
  n1(40 downto 40) &
  n1(39 downto 39) &
  n1(38 downto 38) &
  n1(37 downto 37) &
  n1(36 downto 36) &
  n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(44 downto 44) &
  n1(43 downto 43) &
  n1(42 downto 42);
n4 <= s11_1 & s12_1;
n5 <= n1(44 downto 44);
n6 <= n5 & s12_2;
n7 <= i1(47 downto 47) &
  i1(46 downto 46) &
  i1(45 downto 45);
n8 <= s13_1 & n4;
n9 <= i1(47 downto 47);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_5 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_3 is
port (
i1 : in  unsigned(53 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0));
end entity cf_ldpc_3;
architecture rtl of cf_ldpc_3 is
signal n1 : unsigned(50 downto 0);
signal n2 : unsigned(47 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(16 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(16 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(17 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(17 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(15 downto 0);
signal s12_2 : unsigned(15 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_4 is
port (
i1 : in  unsigned(47 downto 0);
o1 : out unsigned(15 downto 0);
o2 : out unsigned(15 downto 0));
end component cf_ldpc_4;
begin
n1 <= i1(50 downto 50) &
  i1(49 downto 49) &
  i1(48 downto 48) &
  i1(47 downto 47) &
  i1(46 downto 46) &
  i1(45 downto 45) &
  i1(44 downto 44) &
  i1(43 downto 43) &
  i1(42 downto 42) &
  i1(41 downto 41) &
  i1(40 downto 40) &
  i1(39 downto 39) &
  i1(38 downto 38) &
  i1(37 downto 37) &
  i1(36 downto 36) &
  i1(35 downto 35) &
  i1(34 downto 34) &
  i1(33 downto 33) &
  i1(32 downto 32) &
  i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(47 downto 47) &
  n1(46 downto 46) &
  n1(45 downto 45) &
  n1(44 downto 44) &
  n1(43 downto 43) &
  n1(42 downto 42) &
  n1(41 downto 41) &
  n1(40 downto 40) &
  n1(39 downto 39) &
  n1(38 downto 38) &
  n1(37 downto 37) &
  n1(36 downto 36) &
  n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(50 downto 50) &
  n1(49 downto 49) &
  n1(48 downto 48);
n4 <= s11_1 & s12_1;
n5 <= n1(50 downto 50);
n6 <= n5 & s12_2;
n7 <= i1(53 downto 53) &
  i1(52 downto 52) &
  i1(51 downto 51);
n8 <= s13_1 & n4;
n9 <= i1(53 downto 53);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_4 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_2 is
port (
i1 : in  unsigned(59 downto 0);
o1 : out unsigned(19 downto 0);
o2 : out unsigned(19 downto 0));
end entity cf_ldpc_2;
architecture rtl of cf_ldpc_2 is
signal n1 : unsigned(56 downto 0);
signal n2 : unsigned(53 downto 0);
signal n3 : unsigned(2 downto 0);
signal n4 : unsigned(18 downto 0);
signal n5 : unsigned(0 downto 0);
signal n6 : unsigned(18 downto 0);
signal n7 : unsigned(2 downto 0);
signal n8 : unsigned(19 downto 0);
signal n9 : unsigned(0 downto 0);
signal n10 : unsigned(19 downto 0);
signal s11_1 : unsigned(0 downto 0);
signal s12_1 : unsigned(17 downto 0);
signal s12_2 : unsigned(17 downto 0);
signal s13_1 : unsigned(0 downto 0);
component cf_ldpc_12 is
port (
i1 : in  unsigned(2 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_12;
component cf_ldpc_3 is
port (
i1 : in  unsigned(53 downto 0);
o1 : out unsigned(17 downto 0);
o2 : out unsigned(17 downto 0));
end component cf_ldpc_3;
begin
n1 <= i1(56 downto 56) &
  i1(55 downto 55) &
  i1(54 downto 54) &
  i1(53 downto 53) &
  i1(52 downto 52) &
  i1(51 downto 51) &
  i1(50 downto 50) &
  i1(49 downto 49) &
  i1(48 downto 48) &
  i1(47 downto 47) &
  i1(46 downto 46) &
  i1(45 downto 45) &
  i1(44 downto 44) &
  i1(43 downto 43) &
  i1(42 downto 42) &
  i1(41 downto 41) &
  i1(40 downto 40) &
  i1(39 downto 39) &
  i1(38 downto 38) &
  i1(37 downto 37) &
  i1(36 downto 36) &
  i1(35 downto 35) &
  i1(34 downto 34) &
  i1(33 downto 33) &
  i1(32 downto 32) &
  i1(31 downto 31) &
  i1(30 downto 30) &
  i1(29 downto 29) &
  i1(28 downto 28) &
  i1(27 downto 27) &
  i1(26 downto 26) &
  i1(25 downto 25) &
  i1(24 downto 24) &
  i1(23 downto 23) &
  i1(22 downto 22) &
  i1(21 downto 21) &
  i1(20 downto 20) &
  i1(19 downto 19) &
  i1(18 downto 18) &
  i1(17 downto 17) &
  i1(16 downto 16) &
  i1(15 downto 15) &
  i1(14 downto 14) &
  i1(13 downto 13) &
  i1(12 downto 12) &
  i1(11 downto 11) &
  i1(10 downto 10) &
  i1(9 downto 9) &
  i1(8 downto 8) &
  i1(7 downto 7) &
  i1(6 downto 6) &
  i1(5 downto 5) &
  i1(4 downto 4) &
  i1(3 downto 3) &
  i1(2 downto 2) &
  i1(1 downto 1) &
  i1(0 downto 0);
n2 <= n1(53 downto 53) &
  n1(52 downto 52) &
  n1(51 downto 51) &
  n1(50 downto 50) &
  n1(49 downto 49) &
  n1(48 downto 48) &
  n1(47 downto 47) &
  n1(46 downto 46) &
  n1(45 downto 45) &
  n1(44 downto 44) &
  n1(43 downto 43) &
  n1(42 downto 42) &
  n1(41 downto 41) &
  n1(40 downto 40) &
  n1(39 downto 39) &
  n1(38 downto 38) &
  n1(37 downto 37) &
  n1(36 downto 36) &
  n1(35 downto 35) &
  n1(34 downto 34) &
  n1(33 downto 33) &
  n1(32 downto 32) &
  n1(31 downto 31) &
  n1(30 downto 30) &
  n1(29 downto 29) &
  n1(28 downto 28) &
  n1(27 downto 27) &
  n1(26 downto 26) &
  n1(25 downto 25) &
  n1(24 downto 24) &
  n1(23 downto 23) &
  n1(22 downto 22) &
  n1(21 downto 21) &
  n1(20 downto 20) &
  n1(19 downto 19) &
  n1(18 downto 18) &
  n1(17 downto 17) &
  n1(16 downto 16) &
  n1(15 downto 15) &
  n1(14 downto 14) &
  n1(13 downto 13) &
  n1(12 downto 12) &
  n1(11 downto 11) &
  n1(10 downto 10) &
  n1(9 downto 9) &
  n1(8 downto 8) &
  n1(7 downto 7) &
  n1(6 downto 6) &
  n1(5 downto 5) &
  n1(4 downto 4) &
  n1(3 downto 3) &
  n1(2 downto 2) &
  n1(1 downto 1) &
  n1(0 downto 0);
n3 <= n1(56 downto 56) &
  n1(55 downto 55) &
  n1(54 downto 54);
n4 <= s11_1 & s12_1;
n5 <= n1(56 downto 56);
n6 <= n5 & s12_2;
n7 <= i1(59 downto 59) &
  i1(58 downto 58) &
  i1(57 downto 57);
n8 <= s13_1 & n4;
n9 <= i1(59 downto 59);
n10 <= n9 & n6;
s11 : cf_ldpc_12 port map (n3, s11_1);
s12 : cf_ldpc_3 port map (n2, s12_1, s12_2);
s13 : cf_ldpc_12 port map (n7, s13_1);
o2 <= n10;
o1 <= n8;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(19 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(19 downto 0));
end entity cf_ldpc_1;
architecture rtl of cf_ldpc_1 is
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(0 downto 0);
signal n3 : unsigned(19 downto 0) := "00000000000000000000";
signal n4 : unsigned(19 downto 0);
signal n5 : unsigned(19 downto 0) := "00000000000000000000";
signal s6_1 : unsigned(19 downto 0);
signal s7_1 : unsigned(59 downto 0);
signal s8_1 : unsigned(0 downto 0);
signal s9_1 : unsigned(19 downto 0);
signal s9_2 : unsigned(19 downto 0);
component cf_ldpc_85 is
port (
i1 : in  unsigned(19 downto 0);
i2 : in  unsigned(19 downto 0);
i3 : in  unsigned(19 downto 0);
o1 : out unsigned(19 downto 0));
end component cf_ldpc_85;
component cf_ldpc_25 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(59 downto 0));
end component cf_ldpc_25;
component cf_ldpc_14 is
port (
i1 : in  unsigned(19 downto 0);
o1 : out unsigned(0 downto 0));
end component cf_ldpc_14;
component cf_ldpc_2 is
port (
i1 : in  unsigned(59 downto 0);
o1 : out unsigned(19 downto 0);
o2 : out unsigned(19 downto 0));
end component cf_ldpc_2;
begin
n1 <= "1";
n2 <= "0";
process (clock_c) begin
  if rising_edge(clock_c) then
    if n2 = "1" then
      n3 <= "00000000000000000000";
    elsif i1 = "1" then
      n3 <= i2;
    end if;
  end if;
end process;
n4 <= i2 when i1 = "1" else s6_1;
process (clock_c) begin
  if rising_edge(clock_c) then
    if n2 = "1" then
      n5 <= "00000000000000000000";
    elsif n1 = "1" then
      n5 <= n4;
    end if;
  end if;
end process;
s6 : cf_ldpc_85 port map (n3, s9_1, s9_2, s6_1);
s7 : cf_ldpc_25 port map (n5, s7_1);
s8 : cf_ldpc_14 port map (n5, s8_1);
s9 : cf_ldpc_2 port map (s7_1, s9_1, s9_2);
o2 <= n5;
o1 <= s8_1;
end architecture rtl;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity cf_ldpc is
port(
signal clock_c : in std_logic;
signal start_i : in unsigned(0 downto 0);
signal message_i : in unsigned(19 downto 0);
signal valid_o : out unsigned(0 downto 0);
signal message_o : out unsigned(19 downto 0));
end entity cf_ldpc;
architecture rtl of cf_ldpc is
component cf_ldpc_1 is
port (
clock_c : in std_logic;
i1 : in  unsigned(0 downto 0);
i2 : in  unsigned(19 downto 0);
o1 : out unsigned(0 downto 0);
o2 : out unsigned(19 downto 0));
end component cf_ldpc_1;
signal n1 : unsigned(0 downto 0);
signal n2 : unsigned(19 downto 0);
begin
s1 : cf_ldpc_1 port map (clock_c, start_i, message_i, n1, n2);
valid_o <= n1;
message_o <= n2;
end architecture rtl;


